library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity SampleMemory is
	Port ( Clk : in  STD_LOGIC;
	       Write_Enable : in  STD_LOGIC;
	       Write_Addr : in  STD_LOGIC_VECTOR (9 downto 0);
	       Write_Data : in  STD_LOGIC_VECTOR (8 downto 0);
	       Read_Addr : in  STD_LOGIC_VECTOR (9 downto 0);
	       Read_Data : out  STD_LOGIC_VECTOR (8 downto 0) );
end SampleMemory;

architecture Behavioral of SampleMemory is
	Type storage_type is array (0 to 799) of std_logic_vector (8 downto 0);
	Signal samples : storage_type := ("000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000",
	                                  "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000", "000000000");
begin
	
	Read_write : process (Clk)
	begin
		if ( rising_edge(Clk) ) then
			if (Write_Enable = '1') then
				samples(to_integer(unsigned((Write_Addr)))) <= Write_Data;
			end if;
			Read_Data <= samples(to_integer(unsigned((Read_Addr))));
		end if;
	end process;
	
end Behavioral;
